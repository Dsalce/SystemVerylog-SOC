`timescale 1ns / 1ps

package definitions;

import uvm_pkg::*;

`include "uvm_macros.svh"
`include "transaction.sv"
`include "sequencer.sv"
`include "sequence.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include "test.sv"



endpackage : definitions