

class transaction;

  //Declaracion de los datos randomizados
  rand bit  [7:0] A;//data
  rand bit  [7:0] B;//data
  rand bit  [2:0] op;//op
  bit start;
  bit done;
  bit [15:0] result;







endclass
