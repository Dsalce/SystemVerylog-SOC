

package agent;


`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"

 endpackage : agent
